// SPDX-License-Identifier: BSD-3-Clause

(* techmap_celltype = "$_DLATCH_P_" *)
module _80_FET_dlatch_p (CLK, D, Q);
	input  CLK;
	input  D;
	output Q;

endmodule

(* techmap_celltype = "$_DLATCH_N_" *)
module _80_FET_dlatch_n (CLK, D, Q);
	input  CLK;
	input  D;
	output Q;

endmodule


(* techmap_celltype = "$_DFF_N_" *)
module _80_FET_dff_n (CLK, D, Q);
	input  CLK;
	input  D;
	output Q;


endmodule

(* techmap_celltype = "$_DFF_P_" *)
module _80_FET_dff_p (CLK, D, Q);
	input  CLK;
	input  D;
	output Q;

endmodule
