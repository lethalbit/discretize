// SPDX-License-Identifier: BSD-3-Clause

(* techmap_celltype = "$_DFF_N_" *)
module _80_FET_dff_n (C, D, Q, Qn);


endmodule

(* techmap_celltype = "$_DFF_P_" *)
module _80_FET_dff_p (C, D, Q, Qn);


endmodule
